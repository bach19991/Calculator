library ieee;
use ieee.std_logic_1164.all;

entity shiftleft48bit is
port (	a	:	in	std_logic_vector(23 downto 0);
		s	:	in	std_logic_vector(5 downto 0);
		y	:	out	std_logic_vector(47 downto 0));
end shiftleft48bit;

architecture struc of shiftleft48bit is
component mux48to1 is
port(	a0,a1,a2,a3,a4,a5,a6,a7,a8,a9	:	in	std_logic;
		a10,a11,a12,a13,a14,a15,a16		:	in	std_logic;
		a17,a18,a19,a20,a21,a22,a23,a24	:	in	std_logic;
		a25,a26,a27,a28,a29,a30,a31,a32	:	in	std_logic;
		a33,a34,a35,a36,a37,a38,a39,a40	:	in	std_logic;
		a41,a42,a43,a44,a45,a46,a47		:	in	std_logic;
		s0,s1,s2,s3,s4,s5				:	in	std_logic;
		y								:	out	std_logic);
end component;

begin

																																																																				
mux0	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(47));
mux1	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(46));
mux2	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(45));
mux3	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(44));
mux4	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(43));
mux5	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(42));
mux6	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(41));
mux7	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(40));
mux8	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(39));
mux9	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(38));
mux10	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(37));
mux11	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(36));
mux12	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(35));
mux13	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(34));
mux14	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(33));
mux15	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(32));
mux16	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(31));
mux17	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(30));
mux18	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(29));
mux19	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(28));
mux20	: mux48to1 port map('0'  ,'0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(27));
mux21	: mux48to1 port map('0'  ,'0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(26));
mux22	: mux48to1 port map('0'  ,'0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(25));
mux23	: mux48to1 port map('0'  ,a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(24));
mux24	: mux48to1 port map(a(23),a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(23));
mux25	: mux48to1 port map(a(22),a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(22));
mux26	: mux48to1 port map(a(21),a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(21));
mux27	: mux48to1 port map(a(20),a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(20));
mux28	: mux48to1 port map(a(19),a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(19));
mux29	: mux48to1 port map(a(18),a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(18));
mux30	: mux48to1 port map(a(17),a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(17));
mux31	: mux48to1 port map(a(16),a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(16));
mux32	: mux48to1 port map(a(15),a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(15));
mux33	: mux48to1 port map(a(14),a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(14));
mux34	: mux48to1 port map(a(13),a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(13));
mux35	: mux48to1 port map(a(12),a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(12));
mux36	: mux48to1 port map(a(11),a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(11));
mux37	: mux48to1 port map(a(10),a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(10));
mux38	: mux48to1 port map(a(9 ),a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(9 ));
mux39	: mux48to1 port map(a(8 ),a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(8 ));
mux40	: mux48to1 port map(a(7 ),a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(7 ));
mux41	: mux48to1 port map(a(6 ),a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(6 ));
mux42	: mux48to1 port map(a(5 ),a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(5 ));
mux43	: mux48to1 port map(a(4 ),a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(4 ));
mux44	: mux48to1 port map(a(3 ),a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(3 ));
mux45	: mux48to1 port map(a(2 ),a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(2 ));
mux46	: mux48to1 port map(a(1 ),a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(1 ));
mux47	: mux48to1 port map(a(0 ),'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,'0'  ,s(0 ),s(1 ),s(2 ),s(3 ),s(4 ),s(5 ),y(0 ));
																																																										
																																																			
																																										


end struc;

